module testbench_cfc;

endmodule
