module testbench_cfc;
//comment
endmodule
