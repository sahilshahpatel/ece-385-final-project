module testbench_nfc 

endmodule
