module testbench_cfc;
//comment2
endmodule
